module ks_vandana_fp_div_tb();
reg [31:0]a1,b1;
reg clk;
wire [31:0]c1;

ks_vandana_fp_div DUT(a1,b1,c1,clk);
initial begin
$dumpfile("ks_vandana_fp_div.vcd");
$dumpvars(0,ks_vandana_fp_div_tb);
end
initial clk=0;
always #5 clk=~clk;
initial begin
a1=32'b01000010111101111011001100110011;//123.85
b1=32'b01000010001101100000000000000000;//45.5
//123.85/45.5 = 2.721978022
#50
a1=32'b01000010000101110101000011100101;//37.829
b1=32'b01000000000010001110010101100000;//2.139
//37.829/2.139 = 17.68536699
#50
a1=32'b01000010100001101101001101110101;//67.413
b1=32'b01000001000011110001001001101111;//8.942
//67.413/8.942 = 7.538917468
#250 $finish;
end
endmodule
